module LUT_S(addr, out);
	input [5:0] addr;
	output reg [31:0] out;
	always @(addr)
		case(addr)
			6'd0 : out = 5'd7; 
			6'd1 : out = 5'd12;
			6'd2 : out = 5'd17;
			6'd3 : out = 5'd22;
			6'd4 : out = 5'd7; 
			6'd5 : out = 5'd12;
			6'd6 : out = 5'd17;
			6'd7 : out = 5'd22;
			6'd8 : out = 5'd7; 
			6'd9 : out = 5'd12;
			6'd10 : out = 5'd17;
			6'd11 : out = 5'd22;
			6'd12 : out = 5'd7;
			6'd13 : out = 5'd12;
			6'd14 : out = 5'd17;
			6'd15 : out = 5'd22;
			6'd16 : out = 5'd5;
			6'd17 : out = 5'd9;
			6'd18 : out = 5'd14;
			6'd19 : out = 5'd20;
			6'd20 : out = 5'd5;
			6'd21 : out = 5'd9;
			6'd22 : out = 5'd14;
			6'd23 : out = 5'd20;
			6'd14 : out = 5'd5;
			6'd25 : out = 5'd9;
			6'd26 : out = 5'd14;
			6'd27 : out = 5'd20;
			6'd28 : out = 5'd5;
			6'd29 : out = 5'd9;
			6'd30 : out = 5'd14;
			6'd31 : out = 5'd20;
			6'd32 : out = 5'd4;
			6'd33 : out = 5'd11;
			6'd34 : out = 5'd16;
			6'd35 : out = 5'd23;
			6'd36 : out = 5'd4;
			6'd37 : out = 5'd11;
			6'd38 : out = 5'd16;
			6'd39 : out = 5'd23;
			6'd40 : out = 5'd4;
			6'd41 : out = 5'd11;
			6'd42 : out = 5'd16;
			6'd43 : out = 5'd23;
			6'd44 : out = 5'd4;
			6'd45 : out = 5'd11;
			6'd46 : out = 5'd16;
			6'd47 : out = 5'd23;
			6'd48 : out = 5'd6;
			6'd49 : out = 5'd10;
			6'd50 : out = 5'd15;
			6'd51 : out = 5'd21;
			6'd52 : out = 5'd6;
			6'd53 : out = 5'd10;
			6'd54 : out = 5'd15;
			6'd55 : out = 5'd21;
			6'd56 : out = 5'd6;
			6'd57 : out = 5'd10;
			6'd58 : out = 5'd15;
			6'd59 : out = 5'd21;
			6'd60 : out = 5'd6;
			6'd61 : out = 5'd10;
			6'd62 : out = 5'd15;
			6'd63 : out = 5'd21;
	endcase
endmodule

